Library IEEE;
use IEEE.std_logic_1164.all;
Library work;
use work.InstructionSet_12.all;

package rom_program is

  constant pgmadd_w: integer := 10;

  type program_memory_t is array (natural range 0 to 2**pgmadd_w-1) of std_logic_vector(inst_w-1 downto 0);
  constant program : program_memory_t := (
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF",
  X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF"
  ) ;
end package;
